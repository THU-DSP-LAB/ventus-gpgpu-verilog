/*
 * Copyright (c) 2023-2024 C*Core Technology Co.,Ltd,Suzhou.
 * Ventus-RTL is licensed under Mulan PSL v2.
 * You can use this software according to the terms and conditions of the Mulan PSL v2.
 * You may obtain a copy of Mulan PSL v2 at:
 *          http://license.coscl.org.cn/MulanPSL2
 * THIS SOFTWARE IS PROVIDED ON AN "AS IS" BASIS, WITHOUT WARRANTIES OF ANY KIND,
 * EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO NON-INFRINGEMENT,
 * MERCHANTABILITY OR FIT FOR A PARTICULAR PURPOSE.
 * See the Mulan PSL v2 for more details. */
// Author: Zhang, Qi
// Description:
`timescale 1ns/1ns

`include "define.v"

module warp_scheduler (
  input                                     clk                                    ,
  input                                     rst_n                                  ,
                  
  input                                     warpReq_valid_i                        , 
  input      [`TAG_WIDTH-1:0]               warpReq_dispatch2cu_wf_tag_dispatch_i  , //tag of the workgroup
  //input      [`WF_COUNT_WIDTH-1:0]          warpReq_dispatch2cu_wg_wf_count_i      , //sum of warp in a workgroup
  input      [`DEPTH_WARP-1:0]              warpReq_wid_i                          , //warp id
  input      [`MEM_ADDR_WIDTH-1:0]          warpReq_dispatch2cu_start_pc_dispatch_i, //the start pc
                
  input                                     warpRsp_ready_i                        ,
  output                                    warpRsp_valid_o                        , 
  output     [`DEPTH_WARP-1:0]              warpRsp_wid_o                          , //the id of the warp that have ended execution
               
  output     [`DEPTH_WARP-1:0]              wg_id_lookup_o                         , //wid
  input      [`TAG_WIDTH-1:0]               wg_id_tag_i                            , //workgroup's tag
  
  //input                                     pc_req_ready_i                         , 
  output reg                                pc_req_valid_o                         , 
  output     [31:0]                         pc_req_addr_o                          , //fetch pc
  output     [`NUM_FETCH-1:0]               pc_req_mask_o                          ,  
  output     [`DEPTH_WARP-1:0]              pc_req_wid_o                           , //fetch warp id
 
  input                                     pc_rsp_valid_i                         , 
  input      [31:0]                         pc_rsp_addr_i                          , 
  input      [`NUM_FETCH-1:0]               pc_rsp_mask_i                          , 
  input      [`DEPTH_WARP-1:0]              pc_rsp_wid_i                           ,
  input                                     pc_rsp_status_i                        , 

  output                                    branch_ready_o                         , 
  input                                     branch_valid_i                         ,
  input      [`DEPTH_WARP-1:0]              branch_wid_i                           , 
  input                                     branch_jump_i                          , 
  input      [31:0]                         branch_new_pc_i                        , //the pc generated by the branch

  output                                    warp_control_ready_o                   ,
  input                                     warp_control_valid_i                   ,
  input                                     warp_control_simt_stack_op_i           ,
  input      [`DEPTH_WARP-1:0]              warp_control_wid_i                     ,

  input      [`NUM_WARP-1:0]                scoreboard_busy_i                      , 
  //input      [`DEPTH_IBUFFER*`NUM_WARP-1:0] ibuffer_ready_i                        ,
  input      [`NUM_WARP-1:0]                ibuffer_ready_i                        ,
  output     [`NUM_WARP-1:0]                warp_ready_o                           ,

  output                                    flush_valid_o                          , //when branch or warp end, barrier not do this
  output     [`DEPTH_WARP-1:0]              flush_wid_o                            , 

  output                                    flushCache_valid_o                     , //when ibuffer full or icache miss
  output     [`DEPTH_WARP-1:0]              flushCache_wid_o                                   
  );

  wire warp_control_fire;
  wire branch_fire;
  wire warpReq_fire;
  wire warpRsp_fire;
  wire barrier_end;

  wire warp_end;
  wire [`DEPTH_WARP-1:0] warp_end_id;

  wire [`NUM_WARP-1:0] pc_ready;
  reg  [`NUM_WARP-1:0] warp_active;

  wire [31:0]           new_pc_i_tmp  [0:`NUM_WARP-1];
  wire [1:0]            pc_src_i_tmp  [0:`NUM_WARP-1];
  wire [`NUM_FETCH-1:0] mask_i_tmp    [0:`NUM_WARP-1];
  wire [31:0]           pc_next_o_tmp [0:`NUM_WARP-1];
  wire [`NUM_FETCH-1:0] mask_o_tmp    [0:`NUM_WARP-1];

  //reg [`DEPTH_WARP-1:0] current_warp;
  wire [`DEPTH_WARP-1:0] next_warp;

  //reg [`NUM_WARP-1:0] warp_bar_belong [0:`NUM_BLOCK-1]; //active warp
  reg [`NUM_BLOCK*`NUM_WARP-1:0] warp_bar_belong; //[`NUM_WARP-1:0] [0:`NUM_BLOCK-1] active warp
  reg [`NUM_WARP-1:0] warp_bar_data; //barrier

  wire [(`TAG_WIDTH-`WF_COUNT_WIDTH_PER_WG-1):0] new_wg_id,end_wg_id;
  //wire [`WF_COUNT_WIDTH-1:0] new_wg_wf_count; //num of warp in a block

  wire [`NUM_WARP-1:0] next_warp_one_hot;

  wire [`DEPTH_WARP:0] warp_active_tmp;

  //always @(posedge clk or negedge rst_n) begin
  //  if(!rst_n) begin
  //    current_warp <= 'h0;
  //  end
  //  else begin
  //    current_warp <= next_warp;
  //  end
  //end 

  assign branch_ready_o = !flushCache_valid_o;
  assign branch_fire = branch_ready_o && branch_valid_i;

  assign warp_control_ready_o = !branch_fire && !flushCache_valid_o;
  assign warp_control_fire = warp_control_ready_o && warp_control_valid_i;

  assign warp_end = warp_control_fire && warp_control_simt_stack_op_i;
  assign warp_end_id = warp_control_wid_i;

  assign warpReq_fire = warpReq_valid_i;

  assign warpRsp_valid_o = warp_end;
  assign warpRsp_wid_o = warp_end_id;
  assign warpRsp_fire = warpRsp_ready_i && warpRsp_valid_o;

  assign flush_valid_o = (branch_fire && branch_jump_i) || warp_end;
  assign flush_wid_o = (branch_fire && branch_jump_i) ? branch_wid_i : warp_end_id;

  assign flushCache_valid_o = pc_rsp_valid_i && pc_rsp_status_i;
  assign flushCache_wid_o = pc_rsp_wid_i;

  genvar i;
  generate for(i=0;i<`NUM_WARP;i=i+1) begin:B1
    //assign pc_src_i_tmp[i] = ((warpReq_fire && (i == warpReq_wid_i)) || (branch_fire && branch_jump_i && (i == branch_wid_i))) ? 'h1 : 
    //                         ((pc_rsp_valid_i && pc_rsp_status_i && (i == pc_rsp_wid_i)) ? 'h3 :
    //                         ((i == next_warp) ? 'h2 : 'h0));
    assign pc_src_i_tmp[i] = ((warpReq_fire && (i == warpReq_wid_i)) || (branch_fire && branch_jump_i && (i == branch_wid_i))) ? 'h1 : 
                             ((pc_rsp_valid_i && pc_rsp_status_i && (i == pc_rsp_wid_i)) ? 'h3 :
                             ((i == next_warp) ? (((pc_ready=={`NUM_WARP{1'b0}}) && (pc_req_wid_o==next_warp) && (warp_active_tmp > 1)) ? 'h3 :
                             (((pc_ready=={`NUM_WARP{1'b0}}) && (!pc_rsp_valid_i) && (warp_active==1)) ? 'h3 : 'h2)) : 'h0));

    //assign new_pc_i_tmp[i] = (warpReq_fire && (i == warpReq_wid_i)) ? warpReq_dispatch2cu_start_pc_dispatch_i :
    //                         ((pc_rsp_valid_i && pc_rsp_status_i && (i == pc_rsp_wid_i)) ? pc_rsp_addr_i :
    //                         ((branch_fire && branch_jump_i && (i == branch_wid_i)) ? branch_new_pc_i : 'h0));
    assign new_pc_i_tmp[i] = (warpReq_fire && (i == warpReq_wid_i)) ? warpReq_dispatch2cu_start_pc_dispatch_i :
                             ((pc_rsp_valid_i && pc_rsp_status_i && (i == pc_rsp_wid_i)) ? pc_rsp_addr_i :
                             ((branch_fire && branch_jump_i && (i == branch_wid_i)) ? branch_new_pc_i : 
                             (((pc_ready=={`NUM_WARP{1'b0}}) && (i==next_warp) && (pc_req_wid_o==next_warp) && (warp_active_tmp > 1)) ? pc_req_addr_o :
                             (((pc_ready=={`NUM_WARP{1'b0}}) && (!pc_rsp_valid_i) && (warp_active==1)) ? pc_req_addr_o : 'h0))));

    //assign mask_i_tmp[i] = (pc_rsp_valid_i && pc_rsp_status_i && (i == pc_rsp_wid_i)) ? pc_rsp_mask_i : 'h0;
    assign mask_i_tmp[i] = (pc_rsp_valid_i && pc_rsp_status_i && (i == pc_rsp_wid_i)) ? pc_rsp_mask_i : 
                           (((pc_ready=={`NUM_WARP{1'b0}}) && (i==next_warp) && (pc_req_wid_o==next_warp) && (warp_active_tmp > 1)) ? pc_req_mask_o :
                           (((pc_ready=={`NUM_WARP{1'b0}}) && (!pc_rsp_valid_i) && (warp_active==1)) ? pc_req_mask_o : 'h0));

    assign pc_ready[i] = ibuffer_ready_i[i] & warp_active[i];

    pc_control pccontrol(
      .clk      (clk             ),   
      .rst_n    (rst_n           ),  
      .new_pc_i (new_pc_i_tmp[i] ),  
      .pc_src_i (pc_src_i_tmp[i] ),  
      .mask_i   (mask_i_tmp[i]   ),  
      .pc_next_o(pc_next_o_tmp[i]),  
      .mask_o   (mask_o_tmp[i]   )  
      );
  end
  endgenerate 
  
  assign pc_req_addr_o = pc_next_o_tmp[next_warp];
  assign pc_req_wid_o = next_warp;
  assign pc_req_mask_o = mask_o_tmp[next_warp];

  assign wg_id_lookup_o = warp_control_simt_stack_op_i ? warp_end_id : warpRsp_wid_o;
  
  assign new_wg_id=warpReq_dispatch2cu_wf_tag_dispatch_i[`TAG_WIDTH-1:`WF_COUNT_WIDTH_PER_WG];
  //assign new_wg_wf_count=warpReq_dispatch2cu_wg_wf_count_i;
  assign end_wg_id=wg_id_tag_i[`TAG_WIDTH-1:`WF_COUNT_WIDTH_PER_WG];
  
  //genvar j;
  //generate for(j=0;j<`NUM_BLOCK;j=j+1) begin:B2
  //  always @(posedge clk or negedge rst_n) begin
  //    if(!rst_n) begin
  //      warp_bar_belong[j] <= 'h0;
  //    end
  //    else if(warpReq_fire) begin
  //      warp_bar_belong[new_wg_id] <= warp_bar_belong[new_wg_id] | (1 << warpReq_wid_i);
  //    end  
  //    else if(warpRsp_fire) begin
  //      warp_bar_belong[end_wg_id] <= warp_bar_belong[end_wg_id] & (~(1 << warpRsp_wid_o));
  //    end 
  //    else begin
  //      warp_bar_belong[j] <= warp_bar_belong[j];
  //    end 
  //  end 
  //end
  //endgenerate
  //integer j;
  //always @(posedge clk or negedge rst_n) begin
  //    if(!rst_n) begin
  //      for(j=0;j<`NUM_BLOCK;j=j+1) begin:B2
  //        warp_bar_belong[j] <= 'h0;
  //      end 
  //    end
  //    else if(warpReq_fire) begin
  //      warp_bar_belong[new_wg_id] <= warp_bar_belong[new_wg_id] | (1 << warpReq_wid_i);
  //    end  
  //    else if(warpRsp_fire) begin
  //      warp_bar_belong[end_wg_id] <= warp_bar_belong[end_wg_id] & (~(1 << warpRsp_wid_o));
  //    end 
  //    else begin
  //      for(j=0;j<`NUM_BLOCK;j=j+1) begin:B3
  //        warp_bar_belong[j] <= warp_bar_belong[j];
  //      end 
  //    end 
  //end 
  always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
      warp_bar_belong <= 'h0;
    end 
    else if(warpReq_fire) begin
      warp_bar_belong[(`NUM_WARP*(new_wg_id+1)-1) -: `NUM_WARP] <= warp_bar_belong[(`NUM_WARP*(new_wg_id+1)-1) -: `NUM_WARP] | (1<<warpReq_wid_i);
    end 
    else if(warpRsp_fire) begin
      warp_bar_belong[(`NUM_WARP*(end_wg_id+1)-1) -: `NUM_WARP] <= warp_bar_belong[(`NUM_WARP*(end_wg_id+1)-1) -: `NUM_WARP] & (~(1 << warpRsp_wid_o));
    end 
    else begin
      warp_bar_belong <= warp_bar_belong;
    end 
  end 

  assign barrier_end = ((warp_bar_data | (1 << warp_control_wid_i)) == warp_bar_belong[(`NUM_WARP*(end_wg_id+1)-1) -: `NUM_WARP]);

  always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
      warp_bar_data <= 'h0;
    end
    else if(warp_control_fire && (!warp_control_simt_stack_op_i)) begin
      if(!barrier_end) begin
        warp_bar_data <= warp_bar_data | (1 << warp_control_wid_i);
      end 
      else begin
        warp_bar_data <= warp_bar_data & (~warp_bar_belong[(`NUM_WARP*(end_wg_id+1)-1) -: `NUM_WARP]);
      end 
    end
    else begin
      warp_bar_data <= warp_bar_data;
    end
  end 

  always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
      warp_active <= 'h0;
    end 
    else begin
      warp_active <= (warp_active | ((1 << warpReq_wid_i) & {`NUM_WARP{warpReq_fire}})) & (~((1 << warp_end_id) & {`NUM_WARP{warp_end}})); 
    end 
  end

  assign warp_ready_o = (~(warp_bar_data | scoreboard_busy_i | (~warp_active)));


  pop_cnt #(
    .DATA_LEN(`NUM_WARP    ),
    .DATA_WID(`DEPTH_WARP+1)
    ) warp_active_cnt(
    .data_i(warp_active    ),
    .data_o(warp_active_tmp)
    );
  
  //genvar j;
  //generate for(j=0;j<`NUM_WARP;j=j+1) begin:B2
  //  assign pc_ready[j] = ibuffer_ready_i[j] & warp_active[j];
  //end 
  //endgenerate

  fixed_pri_arb #(.ARB_WIDTH(`NUM_WARP)) fixed_arbiter(
    .req  (pc_ready         ),
    .grant(next_warp_one_hot)
    );

  one2bin #(.ONE_WIDTH(`NUM_WARP),.BIN_WIDTH(`DEPTH_WARP)) one_to_bin(
    .oh (next_warp_one_hot),
    .bin(next_warp        )
    );
  
  always @(*) begin
    if(branch_fire && branch_jump_i && (branch_wid_i == next_warp)) begin
      pc_req_valid_o = 1'h0;
    end 
    else begin 
      pc_req_valid_o = pc_ready[next_warp];
    end 
  end 

endmodule
